/*
*Copyright 2020 wy, virusxiewy99@live.cn
*
*ctrl.v - regfile in riscv-5stage cpu
* 
*/

module ctrl (
    input wire clk_i,
    input wire rst_ni
);
    
endmodule