module ex_mem_stage (
    input wire clk,
    input wire rst_ni;
);
    
endmodule