module id_stage (
    input wire clk_i,
    input wire rst_ni,

    input [31:0] instr_i,
    input [31:0] addr,

    output 
);
    
endmodule