module cache (
    ports
);
    
endmodule