module riscv-core (
    input wire clk;
    input wire rst_n;
);
    
endmodule