/*
*Copyright 2020 wy, virusxiewy99@live.cn
*
*csr_regfile.v - csr regfile in riscv-5stage cpu
* 
*/

module csr_regfile (
    input wire clk_;
    input wire rst_ni;
);
    
endmodule