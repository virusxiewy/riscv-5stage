/*
*Copyright 2020 wy, virusxiewy99@live.cn
*
*decoder.v - as the name, it's a simple decoder for RV32I 
* 
*/

module decoder (
    input wire[31:0] instr,

    output wire is_illegal_instr
);
    
endmodule