module riscv_core (
    input wire clk_i;
    input wire rst_ni;
);
    
endmodule