module id_stage (
    input wire clk_i,
    input wire rst_ni;
);
    
endmodule