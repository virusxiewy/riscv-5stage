module frontend (
    input wire clk_i,
    input wire rst_ni,

    input wire 
);
    
endmodule